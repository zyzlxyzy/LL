module chhhh (N1,N5,N9,N12,N15,N18,N23,N26,N29,N32,
N35,N38,N41,N44,N47,N50,N53,N54,N55,N56,
N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,
N69,N70,N73,N74,N75,N76,N77,N78,N79,N80,
N81,N82,N83,N84,N85,N86,N87,N88,N89,N94,
N97,N100,N103,N106,N109,N110,N111,N112,N113,N114,
N115,N118,N121,N124,N127,N130,N133,N134,N135,N138,
N141,N144,N147,N150,N151,N152,N153,N154,N155,N156,
N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,
N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,
N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,
N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,
N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,
N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,
N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,
N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,
N237,N238,N239,N240,N242,N245,N248,N251,N254,N257,
N260,N263,N267,N271,N274,N277,N280,N283,N286,N289,
N293,N296,N299,N303,N307,N310,N313,N316,N319,N322,
N325,N328,N331,N334,N337,N340,N343,N346,N349,N352,
N355,N358,N361,N364,N367,N382,N241_I,N387,N388,N478,
N482,N484,N486,N489,N492,N501,N505,N507,N509,N511,
N513,N515,N517,N519,N535,N537,N539,N541,N543,N545,
N547,N549,N551,N553,N556,N559,N561,N563,N565,N567,
N569,N571,N573,N582,N643,N707,N813,N881,N882,N883,
N884,N885,N889,N945,N1110,N1111,N1112,N1113,N1114,N1489,
N1490,N1781,N10025,N10101,N10102,N10103,N10104,N10109,N10110,N10111,
N10112,N10350,N10351,N10352,N10353,N10574,N10575,N10576,N10628,N10632,
N10641,N10704,N10706,N10711,N10712,N10713,N10714,N10715,N10716,N10717,
N10718,N10729,N10759,N10760,N10761,N10762,N10763,N10827,N10837,N10838,
N10839,N10840,N10868,N10869,N10870,N10871,N10905,N10906,N10907,N10908,
N11333,N11334,N11340,N11342,N241_O,

keybit0,keybit1,keybit2,keybit3,keybit4,keybit5,keybit6,keybit7,keybit8,keybit9,
keybit10,keybit11,keybit12,keybit13,keybit14);


input  N1,N5,N9,N12,N15,N18,N23,N26,N29,N32,
N35,N38,N41,N44,N47,N50,N53,N54,N55,N56,
N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,
N69,N70,N73,N74,N75,N76,N77,N78,N79,N80,
N81,N82,N83,N84,N85,N86,N87,N88,N89,N94,
N97,N100,N103,N106,N109,N110,N111,N112,N113,N114,
N115,N118,N121,N124,N127,N130,N133,N134,N135,N138,
N141,N144,N147,N150,N151,N152,N153,N154,N155,N156,
N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,
N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,
N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,
N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,
N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,
N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,
N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,
N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,
N237,N238,N239,N240,N242,N245,N248,N251,N254,N257,
N260,N263,N267,N271,N274,N277,N280,N283,N286,N289,
N293,N296,N299,N303,N307,N310,N313,N316,N319,N322,
N325,N328,N331,N334,N337,N340,N343,N346,N349,N352,
N355,N358,N361,N364,N367,N382,N241_I,
keybit0,keybit1,keybit2,keybit3,keybit4,keybit5,keybit6,keybit7,keybit8,keybit9,
keybit10,keybit11,keybit12,keybit13,keybit14;


output N387,N388,N478,N482,N484,N486,N489,N492,N501,N505,
N507,N509,N511,N513,N515,N517,N519,N535,N537,N539,
N541,N543,N545,N547,N549,N551,N553,N556,N559,N561,
N563,N565,N567,N569,N571,N573,N582,N643,N707,N813,
N881,N882,N883,N884,N885,N889,N945,N1110,N1111,N1112,
N1113,N1114,N1489,N1490,N1781,N10025,N10101,N10102,N10103,N10104,
N10109,N10110,N10111,N10112,N10350,N10351,N10352,N10353,N10574,N10575,
N10576,N10628,N10632,N10641,N10704,N10706,N10711,N10712,N10713,N10714,
N10715,N10716,N10717,N10718,N10729,N10759,N10760,N10761,N10762,N10763,
N10827,N10837,N10838,N10839,N10840,N10868,N10869,N10870,N10871,N10905,
N10906,N10907,N10908,N11333,N11334,N11340,N11342,N241_O;


wire  N467,N469,N494,N528,N575,N578,N585,N590,N593,N596,
N599,N604,N609,N614,N625,N628,N632,N636,N641,N642,
N644,N651,N657,N660,N666,N672,N673,N674,N676,N682,
N688,N689,N695,N700,N705,N706,N708,N715,N721,N727,
N733,N734,N742,N748,N749,N750,N758,N759,N762,N768,
N774,N780,N786,N794,N800,N806,N812,N814,N821,N827,
N833,N839,N845,N853,N859,N865,N871,N886,N887,N957,
N1028,N1029,N1109,N1115,N1116,N1119,N1125,N1132,N1136,N1141,
N1147,N1154,N1160,N1167,N1174,N1175,N1182,N1189,N1194,N1199,
N1206,N1211,N1218,N1222,N1227,N1233,N1240,N1244,N1249,N1256,
N1263,N1270,N1277,N1284,N1287,N1290,N1293,N1296,N1299,N1302,
N1305,N1308,N1311,N1314,N1317,N1320,N1323,N1326,N1329,N1332,
N1335,N1338,N1341,N1344,N1347,N1350,N1353,N1356,N1359,N1362,
N1365,N1368,N1371,N1374,N1377,N1380,N1383,N1386,N1389,N1392,
N1395,N1398,N1401,N1404,N1407,N1410,N1413,N1416,N1419,N1422,
N1425,N1428,N1431,N1434,N1437,N1440,N1443,N1446,N1449,N1452,
N1455,N1458,N1461,N1464,N1467,N1470,N1473,N1476,N1479,N1482,
N1485,N1537,N1551,N1649,N1703,N1708,N1713,N1721,N1758,N1782,
N1783,N1789,N1793,N1794,N1795,N1796,N1797,N1798,N1799,N1805,
N1811,N1812,N1813,N1814,N1815,N1816,N1817,N1818,N1819,N1820,
N1821,N1822,N1828,N1829,N1830,N1832,N1833,N1834,N1835,N1839,
N1840,N1841,N1842,N1843,N1845,N1851,N1857,N1858,N1859,N1860,
N1861,N1862,N1863,N1864,N1865,N1866,N1867,N1868,N1869,N1870,
N1871,N1872,N1873,N1874,N1875,N1876,N1877,N1878,N1879,N1880,
N1881,N1882,N1883,N1884,N1885,N1892,N1899,N1906,N1913,N1919,
N1926,N1927,N1928,N1929,N1930,N1931,N1932,N1933,N1934,N1935,
N1936,N1937,N1938,N1939,N1940,N1941,N1942,N1943,N1944,N1945,
N1946,N1947,N1953,N1957,N1958,N1959,N1960,N1961,N1962,N1963,
N1965,N1966,N1967,N1968,N1969,N1970,N1971,N1972,N1973,N1974,
N1975,N1976,N1977,N1983,N1989,N1990,N1991,N1992,N1993,N1994,
N1995,N1996,N1997,N2003,N2010,N2011,N2012,N2013,N2014,N2015,
N2016,N2017,N2018,N2019,N2020,N2021,N2022,N2023,N2024,N2031,
N2038,N2045,N2052,N2058,N2064,N2065,N2066,N2067,N2068,N2069,
N2070,N2071,N2072,N2073,N2074,N2081,N2086,N2107,N2108,N2110,
N2111,N2112,N2113,N2114,N2115,N2117,N2171,N2172,N2230,N2231,
N2235,N2239,N2240,N2241,N2242,N2243,N2244,N2245,N2246,N2247,
N2248,N2249,N2250,N2251,N2252,N2253,N2254,N2255,N2256,N2257,
N2267,N2268,N2269,N2274,N2275,N2277,N2278,N2279,N2280,N2281,
N2282,N2283,N2284,N2285,N2286,N2287,N2293,N2299,N2300,N2301,
N2302,N2303,N2304,N2305,N2306,N2307,N2308,N2309,N2315,N2321,
N2322,N2323,N2324,N2325,N2326,N2327,N2328,N2329,N2330,N2331,
N2337,N2338,N2339,N2340,N2341,N2342,N2343,N2344,N2345,N2346,
N2347,N2348,N2349,N2350,N2351,N2352,N2353,N2354,N2355,N2356,
N2357,N2358,N2359,N2360,N2361,N2362,N2363,N2364,N2365,N2366,
N2367,N2368,N2374,N2375,N2376,N2377,N2378,N2379,N2380,N2381,
N2382,N2383,N2384,N2390,N2396,N2397,N2398,N2399,N2400,N2401,
N2402,N2403,N2404,N2405,N2406,N2412,N2418,N2419,N2420,N2421,
N2422,N2423,N2424,N2425,N2426,N2427,N2428,N2429,N2430,N2431,
N2432,N2433,N2434,N2435,N2436,N2437,N2441,N2442,N2446,N2450,
N2454,N2458,N2462,N2466,N2470,N2474,N2478,N2482,N2488,N2496,
N2502,N2508,N2523,N2533,N2537,N2538,N2542,N2546,N2550,N2554,
N2561,N2567,N2573,N2604,N2607,N2611,N2615,N2619,N2626,N2632,
N2638,N2644,N2650,N2653,N2654,N2658,N2662,N2666,N2670,N2674,
N2680,N2688,N2692,N2696,N2700,N2704,N2728,N2729,N2733,N2737,
N2741,N2745,N2749,N2753,N2757,N2761,N2765,N2766,N2769,N2772,
N2775,N2778,N2781,N2784,N2787,N2790,N2793,N2796,N2866,N2867,
N2868,N2869,N2878,N2913,N2914,N2915,N2916,N2917,N2918,N2919,
N2920,N2921,N2922,N2923,N2924,N2925,N2926,N2927,N2928,N2929,
N2930,N2931,N2932,N2933,N2934,N2935,N2936,N2937,N2988,N3005,
N3006,N3007,N3008,N3009,N3020,N3021,N3022,N3023,N3024,N3025,
N3026,N3027,N3028,N3029,N3032,N3033,N3034,N3035,N3036,N3037,
N3038,N3039,N3040,N3041,N3061,N3064,N3067,N3070,N3073,N3080,
N3096,N3097,N3101,N3107,N3114,N3122,N3126,N3130,N3131,N3134,
N3135,N3136,N3137,N3140,N3144,N3149,N3155,N3159,N3167,N3168,
N3169,N3173,N3178,N3184,N3185,N3189,N3195,N3202,N3210,N3211,
N3215,N3221,N3228,N3229,N3232,N3236,N3241,N3247,N3251,N3255,
N3259,N3263,N3267,N3273,N3281,N3287,N3293,N3299,N3303,N3307,
N3311,N3315,N3322,N3328,N3334,N3340,N3343,N3349,N3355,N3361,
N3362,N3363,N3364,N3365,N3366,N3367,N3368,N3369,N3370,N3371,
N3372,N3373,N3374,N3375,N3379,N3380,N3381,N3384,N3390,N3398,
N3404,N3410,N3416,N3420,N3424,N3428,N3432,N3436,N3440,N3444,
N3448,N3452,N3453,N3454,N3458,N3462,N3466,N3470,N3474,N3478,
N3482,N3486,N3487,N3490,N3493,N3496,N3499,N3502,N3507,N3510,
N3515,N3518,N3521,N3524,N3527,N3530,N3535,N3539,N3542,N3545,
N3548,N3551,N3552,N3553,N3557,N3560,N3563,N3566,N3569,N3570,
N3571,N3574,N3577,N3580,N3583,N3586,N3589,N3592,N3595,N3598,
N3601,N3604,N3607,N3610,N3613,N3616,N3619,N3622,N3625,N3628,
N3631,N3634,N3637,N3640,N3643,N3646,N3649,N3652,N3655,N3658,
N3661,N3664,N3667,N3670,N3673,N3676,N3679,N3682,N3685,N3688,
N3691,N3694,N3697,N3700,N3703,N3706,N3709,N3712,N3715,N3718,
N3721,N3724,N3727,N3730,N3733,N3736,N3739,N3742,N3745,N3748,
N3751,N3754,N3757,N3760,N3763,N3766,N3769,N3772,N3775,N3778,
N3781,N3782,N3783,N3786,N3789,N3792,N3795,N3798,N3801,N3804,
N3807,N3810,N3813,N3816,N3819,N3822,N3825,N3828,N3831,N3834,
N3837,N3840,N3843,N3846,N3849,N3852,N3855,N3858,N3861,N3864,
N3867,N3870,N3873,N3876,N3879,N3882,N3885,N3888,N3891,N3953,
N3954,N3955,N3956,N3958,N3964,N4193,N4303,N4308,N4313,N4326,
N4327,N4333,N4334,N4411,N4412,N4463,N4464,N4465,N4466,N4467,
N4468,N4469,N4470,N4471,N4472,N4473,N4474,N4475,N4476,N4477,
N4478,N4479,N4480,N4481,N4482,N4483,N4484,N4485,N4486,N4487,
N4488,N4489,N4490,N4491,N4492,N4493,N4494,N4495,N4496,N4497,
N4498,N4499,N4500,N4501,N4502,N4503,N4504,N4505,N4506,N4507,
N4508,N4509,N4510,N4511,N4512,N4513,N4514,N4515,N4516,N4517,
N4518,N4519,N4520,N4521,N4522,N4523,N4524,N4525,N4526,N4527,
N4528,N4529,N4530,N4531,N4532,N4533,N4534,N4535,N4536,N4537,
N4538,N4539,N4540,N4541,N4542,N4543,N4544,N4545,N4549,N4555,
N4562,N4563,N4566,N4570,N4575,N4576,N4577,N4581,N4586,N4592,
N4593,N4597,N4603,N4610,N4611,N4612,N4613,N4614,N4615,N4616,
N4617,N4618,N4619,N4620,N4621,N4622,N4623,N4624,N4625,N4626,
N4627,N4628,N4629,N4630,N4631,N4632,N4633,N4634,N4635,N4636,
N4637,N4638,N4639,N4640,N4641,N4642,N4643,N4644,N4645,N4646,
N4647,N4648,N4649,N4650,N4651,N4652,N4653,N4656,N4657,N4661,
N4667,N4674,N4675,N4678,N4682,N4687,N4693,N4694,N4695,N4696,
N4697,N4698,N4699,N4700,N4701,N4702,N4706,N4711,N4717,N4718,
N4722,N4728,N4735,N4743,N4744,N4745,N4746,N4747,N4748,N4749,
N4750,N4751,N4752,N4753,N4754,N4755,N4756,N4757,N4758,N4759,
N4760,N4761,N4762,N4763,N4764,N4765,N4766,N4767,N4768,N4769,
N4775,N4776,N4777,N4778,N4779,N4780,N4781,N4782,N4783,N4784,
N4789,N4790,N4793,N4794,N4795,N4796,N4799,N4800,N4801,N4802,
N4803,N4806,N4809,N4810,N4813,N4814,N4817,N4820,N4823,N4826,
N4829,N4832,N4835,N4838,N4841,N4844,N4847,N4850,N4853,N4856,
N4859,N4862,N4865,N4868,N4871,N4874,N4877,N4880,N4883,N4886,
N4889,N4892,N4895,N4898,N4901,N4904,N4907,N4910,N4913,N4916,
N4919,N4922,N4925,N4928,N4931,N4934,N4937,N4940,N4943,N4946,
N4949,N4952,N4955,N4958,N4961,N4964,N4967,N4970,N4973,N4976,
N4979,N4982,N4985,N4988,N4991,N4994,N4997,N5000,N5003,N5006,
N5009,N5012,N5015,N5018,N5021,N5024,N5027,N5030,N5033,N5036,
N5039,N5042,N5045,N5046,N5047,N5048,N5049,N5052,N5055,N5058,
N5061,N5064,N5065,N5066,N5067,N5068,N5071,N5074,N5077,N5080,
N5083,N5086,N5089,N5092,N5095,N5098,N5101,N5104,N5107,N5110,
N5111,N5112,N5113,N5114,N5117,N5120,N5123,N5126,N5129,N5132,
N5135,N5138,N5141,N5144,N5147,N5150,N5153,N5156,N5159,N5162,
N5165,N5166,N5167,N5168,N5169,N5170,N5171,N5172,N5173,N5174,
N5175,N5176,N5177,N5178,N5179,N5180,N5181,N5182,N5183,N5184,
N5185,N5186,N5187,N5188,N5189,N5190,N5191,N5192,N5193,N5196,
N5197,N5198,N5199,N5200,N5201,N5202,N5203,N5204,N5205,N5206,
N5207,N5208,N5209,N5210,N5211,N5212,N5213,N5283,N5284,N5285,
N5286,N5287,N5288,N5289,N5290,N5291,N5292,N5293,N5294,N5295,
N5296,N5297,N5298,N5299,N5300,N5314,N5315,N5316,N5317,N5318,
N5319,N5320,N5321,N5322,N5323,N5324,N5363,N5364,N5365,N5366,
N5367,N5425,N5426,N5427,N5429,N5430,N5431,N5432,N5433,N5451,
N5452,N5453,N5454,N5455,N5456,N5457,N5469,N5474,N5475,N5476,
N5477,N5571,N5572,N5573,N5574,N5584,N5585,N5586,N5587,N5602,
N5603,N5604,N5605,N5631,N5632,N5640,N5654,N5670,N5683,N5690,
N5697,N5707,N5718,N5728,N5735,N5736,N5740,N5744,N5747,N5751,
N5755,N5758,N5762,N5766,N5769,N5770,N5771,N5778,N5789,N5799,
N5807,N5821,N5837,N5850,N5856,N5863,N5870,N5881,N5892,N5898,
N5905,N5915,N5926,N5936,N5943,N5944,N5945,N5946,N5947,N5948,
N5949,N5950,N5951,N5952,N5953,N5954,N5955,N5956,N5957,N5958,
N5959,N5960,N5966,N5967,N5968,N5969,N5970,N5971,N5972,N5973,
N5974,N5975,N5976,N5977,N5978,N5979,N5980,N5981,N5989,N5990,
N5991,N5996,N6000,N6003,N6009,N6014,N6018,N6021,N6022,N6023,
N6024,N6025,N6026,N6027,N6028,N6029,N6030,N6031,N6032,N6033,
N6034,N6035,N6036,N6037,N6038,N6039,N6040,N6041,N6047,N6052,
N6056,N6059,N6060,N6061,N6062,N6063,N6064,N6065,N6066,N6067,
N6068,N6069,N6070,N6071,N6072,N6073,N6074,N6075,N6076,N6077,
N6078,N6079,N6083,N6087,N6090,N6091,N6092,N6093,N6094,N6095,
N6096,N6097,N6098,N6099,N6100,N6101,N6102,N6103,N6104,N6105,
N6106,N6107,N6108,N6109,N6110,N6111,N6112,N6113,N6114,N6115,
N6116,N6117,N6118,N6119,N6120,N6121,N6122,N6123,N6124,N6125,
N6126,N6127,N6131,N6135,N6136,N6137,N6141,N6145,N6148,N6149,
N6150,N6151,N6152,N6153,N6154,N6155,N6156,N6157,N6158,N6159,
N6160,N6161,N6162,N6163,N6164,N6165,N6166,N6170,N6174,N6177,
N6181,N6182,N6183,N6184,N6185,N6186,N6187,N6188,N6189,N6190,
N6191,N6192,N6193,N6194,N6195,N6196,N6199,N6202,N6203,N6204,
N6207,N6210,N6213,N6214,N6217,N6220,N6223,N6224,N6225,N6226,
N6227,N6228,N6229,N6230,N6231,N6232,N6235,N6236,N6239,N6240,
N6241,N6242,N6243,N6246,N6249,N6252,N6255,N6256,N6257,N6258,
N6259,N6260,N6261,N6262,N6263,N6266,N6540,N6541,N6542,N6543,
N6544,N6545,N6546,N6547,N6555,N6556,N6557,N6558,N6559,N6560,
N6561,N6569,N6594,N6595,N6596,N6597,N6598,N6599,N6600,N6601,
N6602,N6603,N6604,N6605,N6606,N6621,N6622,N6623,N6624,N6625,
N6626,N6627,N6628,N6629,N6639,N6640,N6641,N6642,N6643,N6644,
N6645,N6646,N6647,N6648,N6649,N6650,N6651,N6652,N6653,N6654,
N6655,N6656,N6657,N6658,N6659,N6660,N6661,N6668,N6677,N6678,
N6679,N6680,N6681,N6682,N6683,N6684,N6685,N6686,N6687,N6688,
N6689,N6690,N6702,N6703,N6704,N6705,N6706,N6707,N6708,N6709,
N6710,N6711,N6712,N6729,N6730,N6731,N6732,N6733,N6734,N6735,
N6736,N6741,N6742,N6743,N6744,N6751,N6752,N6753,N6754,N6755,
N6756,N6757,N6758,N6761,N6762,N6766,N6767,N6768,N6769,N6770,
N6771,N6772,N6773,N6774,N6775,N6776,N6777,N6778,N6779,N6780,
N6781,N6782,N6783,N6784,N6787,N6788,N6789,N6790,N6791,N6792,
N6793,N6794,N6795,N6796,N6797,N6800,N6803,N6806,N6809,N6812,
N6815,N6818,N6821,N6824,N6827,N6830,N6833,N6836,N6837,N6838,
N6839,N6840,N6841,N6842,N6843,N6844,N6845,N6848,N6849,N6850,
N6851,N6852,N6853,N6854,N6855,N6856,N6857,N6858,N6859,N6860,
N6861,N6862,N6863,N6864,N6865,N6866,N6867,N6870,N6871,N6872,
N6873,N6874,N6875,N6876,N6877,N6878,N6879,N6880,N6881,N6884,
N6885,N6886,N6887,N6888,N6889,N6890,N6891,N6892,N6893,N6894,
N6901,N6912,N6923,N6929,N6936,N6946,N6957,N6967,N6968,N6969,
N6970,N6977,N6988,N6998,N7006,N7020,N7036,N7049,N7055,N7056,
N7057,N7060,N7061,N7062,N7063,N7064,N7065,N7066,N7067,N7068,
N7073,N7077,N7080,N7086,N7091,N7095,N7098,N7099,N7100,N7103,
N7104,N7105,N7106,N7107,N7114,N7125,N7136,N7142,N7149,N7159,
N7170,N7180,N7187,N7188,N7191,N7194,N7198,N7202,N7205,N7209,
N7213,N7216,N7219,N7222,N7229,N7240,N7250,N7258,N7272,N7288,
N7301,N7307,N7314,N7318,N7322,N7325,N7328,N7331,N7334,N7337,
N7340,N7343,N7346,N7351,N7355,N7358,N7364,N7369,N7373,N7376,
N7377,N7378,N7381,N7384,N7387,N7391,N7394,N7398,N7402,N7405,
N7408,N7411,N7414,N7417,N7420,N7423,N7426,N7429,N7432,N7435,
N7438,N7441,N7444,N7447,N7450,N7453,N7456,N7459,N7462,N7465,
N7468,N7471,N7474,N7477,N7478,N7479,N7482,N7485,N7488,N7491,
N7494,N7497,N7500,N7503,N7506,N7509,N7512,N7515,N7518,N7521,
N7524,N7527,N7530,N7533,N7536,N7539,N7542,N7545,N7548,N7551,
N7552,N7553,N7556,N7557,N7558,N7559,N7560,N7563,N7566,N7569,
N7572,N7573,N7574,N7577,N7580,N7581,N7582,N7585,N7588,N7591,
N7609,N7613,N7620,N7649,N7650,N7655,N7659,N7668,N7671,N7744,
N7822,N7825,N7826,N7852,N8114,N8117,N8131,N8134,N8144,N8145,
N8146,N8156,N8166,N8169,N8183,N8186,N8196,N8200,N8204,N8208,
N8216,N8217,N8218,N8219,N8232,N8233,N8242,N8243,N8244,N8245,
N8246,N8247,N8248,N8249,N8250,N8251,N8252,N8253,N8254,N8260,
N8261,N8262,N8269,N8274,N8275,N8276,N8277,N8278,N8279,N8280,
N8281,N8282,N8283,N8284,N8285,N8288,N8294,N8295,N8296,N8297,
N8298,N8307,N8315,N8317,N8319,N8321,N8322,N8323,N8324,N8325,
N8326,N8333,N8337,N8338,N8339,N8340,N8341,N8342,N8343,N8344,
N8345,N8346,N8347,N8348,N8349,N8350,N8351,N8352,N8353,N8354,
N8355,N8356,N8357,N8358,N8365,N8369,N8370,N8371,N8372,N8373,
N8374,N8375,N8376,N8377,N8378,N8379,N8380,N8381,N8382,N8383,
N8384,N8385,N8386,N8387,N8388,N8389,N8390,N8391,N8392,N8393,
N8394,N8404,N8405,N8409,N8410,N8411,N8412,N8415,N8416,N8417,
N8418,N8421,N8430,N8433,N8434,N8435,N8436,N8437,N8438,N8439,
N8440,N8441,N8442,N8443,N8444,N8447,N8448,N8449,N8450,N8451,
N8452,N8453,N8454,N8455,N8456,N8457,N8460,N8463,N8466,N8469,
N8470,N8471,N8474,N8477,N8480,N8483,N8484,N8485,N8488,N8489,
N8490,N8491,N8492,N8493,N8494,N8495,N8496,N8497,N8500,N8501,
N8502,N8503,N8504,N8505,N8506,N8507,N8508,N8509,N8510,N8511,
N8512,N8513,N8514,N8515,N8516,N8517,N8518,N8519,N8522,N8525,
N8528,N8531,N8534,N8537,N8538,N8539,N8540,N8541,N8545,N8546,
N8547,N8548,N8551,N8552,N8553,N8554,N8555,N8558,N8561,N8564,
N8565,N8566,N8569,N8572,N8575,N8578,N8579,N8580,N8583,N8586,
N8589,N8592,N8595,N8598,N8601,N8604,N8607,N8608,N8609,N8610,
N8615,N8616,N8617,N8618,N8619,N8624,N8625,N8626,N8627,N8632,
N8633,N8634,N8637,N8638,N8639,N8644,N8645,N8646,N8647,N8648,
N8653,N8654,N8655,N8660,N8663,N8666,N8669,N8672,N8675,N8678,
N8681,N8684,N8687,N8690,N8693,N8696,N8699,N8702,N8705,N8708,
N8711,N8714,N8717,N8718,N8721,N8724,N8727,N8730,N8733,N8734,
N8735,N8738,N8741,N8744,N8747,N8750,N8753,N8754,N8755,N8756,
N8757,N8760,N8763,N8766,N8769,N8772,N8775,N8778,N8781,N8784,
N8787,N8790,N8793,N8796,N8799,N8802,N8805,N8808,N8811,N8814,
N8815,N8816,N8817,N8818,N8840,N8857,N8861,N8862,N8863,N8864,
N8865,N8866,N8871,N8874,N8878,N8879,N8880,N8881,N8882,N8883,
N8884,N8885,N8886,N8887,N8888,N8898,N8902,N8920,N8924,N8927,
N8931,N8943,N8950,N8956,N8959,N8960,N8963,N8966,N8991,N8992,
N8995,N8996,N9001,N9005,N9024,N9025,N9029,N9035,N9053,N9054,
N9064,N9065,N9066,N9067,N9068,N9071,N9072,N9073,N9074,N9077,
N9079,N9082,N9083,N9086,N9087,N9088,N9089,N9092,N9093,N9094,
N9095,N9098,N9099,N9103,N9107,N9111,N9117,N9127,N9146,N9149,
N9159,N9160,N9161,N9165,N9169,N9173,N9179,N9180,N9181,N9182,
N9183,N9193,N9203,N9206,N9220,N9223,N9234,N9235,N9236,N9237,
N9238,N9242,N9243,N9244,N9245,N9246,N9247,N9248,N9249,N9250,
N9251,N9252,N9256,N9257,N9258,N9259,N9260,N9261,N9262,N9265,
N9268,N9271,N9272,N9273,N9274,N9275,N9276,N9280,N9285,N9286,
N9287,N9288,N9290,N9292,N9294,N9296,N9297,N9298,N9299,N9300,
N9301,N9307,N9314,N9315,N9318,N9319,N9320,N9321,N9322,N9323,
N9324,N9326,N9332,N9339,N9344,N9352,N9354,N9356,N9358,N9359,
N9360,N9361,N9362,N9363,N9364,N9365,N9366,N9367,N9368,N9369,
N9370,N9371,N9372,N9375,N9381,N9382,N9383,N9384,N9385,N9392,
N9393,N9394,N9395,N9396,N9397,N9398,N9399,N9400,N9401,N9402,
N9407,N9408,N9412,N9413,N9414,N9415,N9416,N9417,N9418,N9419,
N9420,N9421,N9422,N9423,N9426,N9429,N9432,N9435,N9442,N9445,
N9454,N9455,N9456,N9459,N9460,N9461,N9462,N9465,N9466,N9467,
N9468,N9473,N9476,N9477,N9478,N9485,N9488,N9493,N9494,N9495,
N9498,N9499,N9500,N9505,N9506,N9507,N9508,N9509,N9514,N9515,
N9516,N9517,N9520,N9526,N9531,N9539,N9540,N9541,N9543,N9551,
N9555,N9556,N9557,N9560,N9561,N9562,N9563,N9564,N9565,N9566,
N9567,N9568,N9569,N9570,N9571,N9575,N9579,N9581,N9582,N9585,
N9591,N9592,N9593,N9594,N9595,N9596,N9597,N9598,N9599,N9600,
N9601,N9602,N9603,N9604,N9605,N9608,N9611,N9612,N9613,N9614,
N9615,N9616,N9617,N9618,N9621,N9622,N9623,N9624,N9626,N9629,
N9632,N9635,N9642,N9645,N9646,N9649,N9650,N9653,N9656,N9659,
N9660,N9661,N9662,N9663,N9666,N9667,N9670,N9671,N9674,N9675,
N9678,N9679,N9682,N9685,N9690,N9691,N9692,N9695,N9698,N9702,
N9707,N9710,N9711,N9714,N9715,N9716,N9717,N9720,N9721,N9722,
N9723,N9726,N9727,N9732,N9733,N9734,N9735,N9736,N9737,N9738,
N9739,N9740,N9741,N9742,N9754,N9758,N9762,N9763,N9764,N9765,
N9766,N9767,N9768,N9769,N9773,N9774,N9775,N9779,N9784,N9785,
N9786,N9790,N9791,N9795,N9796,N9797,N9798,N9799,N9800,N9801,
N9802,N9803,N9805,N9806,N9809,N9813,N9814,N9815,N9816,N9817,
N9820,N9825,N9826,N9827,N9828,N9829,N9830,N9835,N9836,N9837,
N9838,N9846,N9847,N9862,N9863,N9866,N9873,N9876,N9890,N9891,
N9892,N9893,N9894,N9895,N9896,N9897,N9898,N9899,N9900,N9901,
N9902,N9903,N9904,N9905,N9906,N9907,N9908,N9909,N9910,N9911,
N9917,N9923,N9924,N9925,N9932,N9935,N9938,N9939,N9945,N9946,
N9947,N9948,N9949,N9953,N9954,N9955,N9956,N9957,N9958,N9959,
N9960,N9961,N9964,N9967,N9968,N9969,N9970,N9971,N9972,N9973,
N9974,N9975,N9976,N9977,N9978,N9979,N9982,N9983,N9986,N9989,
N9992,N9995,N9996,N9997,N9998,N9999,N10002,N10003,N10006,N10007,
N10010,N10013,N10014,N10015,N10016,N10017,N10018,N10019,N10020,N10021,
N10022,N10023,N10024,N10026,N10028,N10032,N10033,N10034,N10035,N10036,
N10037,N10038,N10039,N10040,N10041,N10042,N10043,N10050,N10053,N10054,
N10055,N10056,N10057,N10058,N10059,N10060,N10061,N10062,N10067,N10070,
N10073,N10076,N10077,N10082,N10083,N10084,N10085,N10086,N10093,N10094,
N10105,N10106,N10107,N10108,N10113,N10114,N10115,N10116,N10119,N10124,
N10130,N10131,N10132,N10133,N10134,N10135,N10136,N10137,N10138,N10139,
N10140,N10141,N10148,N10155,N10156,N10157,N10158,N10159,N10160,N10161,
N10162,N10163,N10164,N10165,N10170,N10173,N10176,N10177,N10178,N10179,
N10180,N10183,N10186,N10189,N10192,N10195,N10196,N10197,N10200,N10203,
N10204,N10205,N10206,N10212,N10213,N10230,N10231,N10232,N10233,N10234,
N10237,N10238,N10239,N10240,N10241,N10242,N10247,N10248,N10259,N10264,
N10265,N10266,N10267,N10268,N10269,N10270,N10271,N10272,N10273,N10278,
N10279,N10280,N10281,N10282,N10283,N10287,N10288,N10289,N10290,N10291,
N10292,N10293,N10294,N10295,N10296,N10299,N10300,N10301,N10306,N10307,
N10308,N10311,N10314,N10315,N10316,N10317,N10318,N10321,N10324,N10325,
N10326,N10327,N10328,N10329,N10330,N10331,N10332,N10333,N10334,N10337,
N10338,N10339,N10340,N10341,N10344,N10354,N10357,N10360,N10367,N10375,
N10381,N10388,N10391,N10399,N10402,N10406,N10409,N10412,N10415,N10419,
N10422,N10425,N10428,N10431,N10432,N10437,N10438,N10439,N10440,N10441,
N10444,N10445,N10450,N10451,N10455,N10456,N10465,N10466,N10479,N10497,
N10509,N10512,N10515,N10516,N10517,N10518,N10519,N10522,N10525,N10528,
N10531,N10534,N10535,N10536,N10539,N10542,N10543,N10544,N10545,N10546,
N10547,N10548,N10549,N10550,N10551,N10552,N10553,N10554,N10555,N10556,
N10557,N10558,N10559,N10560,N10561,N10562,N10563,N10564,N10565,N10566,
N10567,N10568,N10569,N10570,N10571,N10572,N10573,N10577,N10581,N10582,
N10583,N10587,N10588,N10589,N10594,N10595,N10596,N10597,N10598,N10602,
N10609,N10610,N10621,N10626,N10627,N10629,N10631,N10637,N10638,N10639,
N10640,N10642,N10643,N10644,N10645,N10647,N10648,N10649,N10652,N10659,
N10662,N10665,N10668,N10671,N10672,N10673,N10674,N10675,N10678,N10681,
N10682,N10683,N10684,N10685,N10686,N10687,N10688,N10689,N10690,N10691,
N10694,N10695,N10696,N10697,N10698,N10701,N10705,N10707,N10708,N10709,
N10710,N10719,N10720,N10730,N10731,N10737,N10738,N10739,N10746,N10747,
N10748,N10749,N10750,N10753,N10754,N10764,N10765,N10766,N10767,N10768,
N10769,N10770,N10771,N10772,N10773,N10774,N10775,N10776,N10778,N10781,
N10784,N10789,N10792,N10796,N10797,N10798,N10799,N10800,N10803,N10806,
N10809,N10812,N10815,N10816,N10817,N10820,N10823,N10824,N10825,N10826,
N10832,N10833,N10834,N10835,N10836,N10845,N10846,N10857,N10862,N10863,
N10864,N10865,N10866,N10867,N10872,N10873,N10874,N10875,N10876,N10879,
N10882,N10883,N10884,N10885,N10886,N10887,N10888,N10889,N10890,N10891,
N10892,N10895,N10896,N10897,N10898,N10899,N10902,N10909,N10910,N10915,
N10916,N10917,N10918,N10919,N10922,N10923,N10928,N10931,N10934,N10935,
N10936,N10937,N10938,N10941,N10944,N10947,N10950,N10953,N10954,N10955,
N10958,N10961,N10962,N10963,N10964,N10969,N10970,N10981,N10986,N10987,
N10988,N10989,N10990,N10991,N10992,N10995,N10998,N10999,N11000,N11001,
N11002,N11003,N11004,N11005,N11006,N11007,N11008,N11011,N11012,N11013,
N11014,N11015,N11018,N11023,N11024,N11027,N11028,N11029,N11030,N11031,
N11034,N11035,N11040,N11041,N11042,N11043,N11044,N11047,N11050,N11053,
N11056,N11059,N11062,N11065,N11066,N11067,N11070,N11073,N11074,N11075,
N11076,N11077,N11078,N11095,N11098,N11099,N11100,N11103,N11106,N11107,
N11108,N11109,N11110,N11111,N11112,N11113,N11114,N11115,N11116,N11117,
N11118,N11119,N11120,N11121,N11122,N11123,N11124,N11127,N11130,N11137,
N11138,N11139,N11140,N11141,N11142,N11143,N11144,N11145,N11152,N11153,
N11154,N11155,N11156,N11159,N11162,N11165,N11168,N11171,N11174,N11177,
N11180,N11183,N11184,N11185,N11186,N11187,N11188,N11205,N11210,N11211,
N11212,N11213,N11214,N11215,N11216,N11217,N11218,N11219,N11220,N11222,
N11223,N11224,N11225,N11226,N11227,N11228,N11229,N11231,N11232,N11233,
N11236,N11239,N11242,N11243,N11244,N11245,N11246,N11250,N11252,N11257,
N11260,N11261,N11262,N11263,N11264,N11265,N11267,N11268,N11269,N11270,
N11272,N11277,N11278,N11279,N11280,N11282,N11283,N11284,N11285,N11286,
N11288,N11289,N11290,N11291,N11292,N11293,N11294,N11295,N11296,N11297,
N11298,N11299,N11302,N11307,N11308,N11309,N11312,N11313,N11314,N11315,
N11316,N11317,N11320,N11321,N11323,N11327,N11328,N11329,N11331,N11335,
N11336,N11337,N11338,N11339,N11341,
keypoint0,keypoint1,keypoint2,keypoint3,keypoint4,keypoint5,keypoint6,keypoint7,keypoint8,keypoint9,
keypoint10,keypoint11,keypoint12,keypoint13,keypoint14;


not A (n1, n2);
not B (n1, n3);
not C (n1, n4);

endmodule